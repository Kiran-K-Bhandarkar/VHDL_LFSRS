LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.all;

ENTITY LFSR_TB IS 
END ENTITY LFSR_TB;

ARCHITECTURE BEHAVIORAL OF LFSR_TB IS
SIGNAL CLK, RST, SEED_IN, EN : STD_LOGIC;
SIGNAL LFSR_SEED, OUTPUT     : STD_LOGIC_VECTOR(4 DOWNTO 0);
     
CONSTANT CLK_PERIOD : TIME := 1 NS;

BEGIN
   UUT: ENTITY WORK.LFSR_5BIT
    PORT MAP
      ( CLK       => CLK,
		RST       => RST,
		SEED_IN   => SEED_IN,
		EN        => EN,
		LFSR_SEED => LFSR_SEED,
		OUTPUT    => OUTPUT
	  );
		
  CLK_PROCESS :PROCESS
   BEGIN
        CLK <= '0';
        WAIT FOR CLK_PERIOD/2;  
        CLK <= '1';
        WAIT FOR CLK_PERIOD/2; 
   END PROCESS;
   
   TEST_PROCESS: PROCESS
     BEGIN  
	   RST <= '0';
	   WAIT FOR CLK_PERIOD;
	   RST <= '1';
	   WAIT FOR CLK_PERIOD;
	   SEED_IN <= '1';
	   LFSR_SEED <= "10000";
	   WAIT FOR CLK_PERIOD;
	   SEED_IN <= '0';
	   WAIT FOR CLK_PERIOD;
	   EN <= '1';
	   WAIT;
	   END PROCESS;
END BEHAVIORAL;

